library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity encryptDecrypt8 is
port(
        clk : in std_logic;

        -- specify your own signals
        );
end encryptDecrypt8;

architecture behav of encryptDecrypt8 is

-- Specify Components here..

-- .. End of Component Specify

-- Specify Signals here..

-- EndofSignalSpecification

begin
-- put your own code here ..

-- EndofCode

end behav;