library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
 
entity full_adder is
port (
        a  : in std_logic;
        b  : in std_logic;
        c_in : in std_logic;
        s   : out std_logic;
        c_out : out std_logic);
end full_adder;

architecture behav of full_adder is
 
-- Specify Signals here..

-- EndofSignalSpecification

begin
-- put your own code here ..

-- EndofCode

end behav;